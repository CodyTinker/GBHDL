//--------------------------------------------------------------------------------//
//  Project Name : GB80                                                           //
//  Module Name  : controller_sequencer.v                                          //
//  Create Date  : August, 2016                                                   //
//  Author       : Kevin Millar                                                   //
//                 Cody Tinker                                                    //
//                                                                                //
//  Description:   Processor Controller Sequencer.                                //
//                                                                                //
//  Dependencies:  None                                                           //
//                                                                                //
//--------------------------------------------------------------------------------//
//  Revision 0.01 - File Created                                                  //
//--------------------------------------------------------------------------------//
module controller_sequencer #(
)(
)
