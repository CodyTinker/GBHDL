//--------------------------------------------------------------------------------//
//  Project Name : GB80                                                           //
//  Module Name  : decoder.v                                                      //
//  Create Date  : August, 2016                                                   //
//  Author       : Kevin Millar                                                   //
//                 Cody Tinker                                                    //
//                                                                                //
//  Description:   Processor Decoder module.                                      //
//                                                                                //
//  Dependencies:  None                                                           //
//                                                                                //
//--------------------------------------------------------------------------------//
//  Revision 0.01 - File Created                                                  //
//--------------------------------------------------------------------------------//
module decoder #(
)(
)

endmodule